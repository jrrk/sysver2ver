`timescale 1 ns / 1 ps
// `default_nettype none
// `define DEBUGNETS
// `define DEBUGREGS
// `define DEBUGASM
// `define DEBUG

`ifdef DEBUG
  `define debug(debug_command) debug_command
`else
  `define debug(debug_command)
`endif

`ifdef FORMAL
  `define FORMAL_KEEP (* keep *)
  `define assert(assert_expr) assert(assert_expr)
`else
  `ifdef DEBUGNETS
    `define FORMAL_KEEP (* keep *)
  `else
    `define FORMAL_KEEP
  `endif
  `define assert(assert_expr) empty_statement
`endif

// uncomment this for register file in extra module
// `define PICORV32_REGS picorv32_regs

// this macro can be used to check if the verilog files in your
// design are read in the correct order.
`define PICORV32_V


/***************************************************************
 * picorv32
 ***************************************************************/

module irq #(
	parameter [ 0:0] ENABLE_COUNTERS = 1,
	parameter [ 0:0] ENABLE_COUNTERS64 = 1,
	parameter [ 0:0] ENABLE_REGS_16_31 = 1,
	parameter [ 0:0] ENABLE_REGS_DUALPORT = 1,
	parameter [ 0:0] LATCHED_MEM_RDATA = 0,
	parameter [ 0:0] TWO_STAGE_SHIFT = 1,
	parameter [ 0:0] BARREL_SHIFTER = 0,
	parameter [ 0:0] TWO_CYCLE_COMPARE = 0,
	parameter [ 0:0] TWO_CYCLE_ALU = 0,
	parameter [ 0:0] COMPRESSED_ISA = 1,
	parameter [ 0:0] CATCH_MISALIGN = 1,
	parameter [ 0:0] CATCH_ILLINSN = 1,
	parameter [ 0:0] ENABLE_PCPI = 0,
	parameter [ 0:0] ENABLE_MUL = 1,
	parameter [ 0:0] ENABLE_FAST_MUL = 0,
	parameter [ 0:0] ENABLE_DIV = 1,
	parameter [ 0:0] ENABLE_IRQ = 1,
	parameter [ 0:0] ENABLE_IRQ_QREGS = 1,
	parameter [ 0:0] ENABLE_IRQ_TIMER = 1,
	parameter [ 0:0] ENABLE_TRACE = 1,
	parameter [ 0:0] REGS_INIT_ZERO = 0,
	parameter [31:0] MASKED_IRQ = 32'h 0000_0000,
	parameter [31:0] LATCHED_IRQ = 32'h ffff_ffff,
	parameter [31:0] PROGADDR_RESET = 32'h 0000_0000,
	parameter [31:0] PROGADDR_IRQ = 32'h 0000_0010,
	parameter [31:0] STACKADDR = 32'h ffff_ffff,
	parameter integer regindex_bits = (ENABLE_REGS_16_31 ? 5 : 4) + ENABLE_IRQ*ENABLE_IRQ_QREGS
) (
	input 			       clk, resetn,
	output reg 		       trap,

	input [31:0] 		       mem_rdata,

	// IRQ Interface
	input [31:0] 		       irq,
	output reg [31:0] 	       eoi,

	// Trace Interface
   	input 			       decoder_trigger,
	input 			       do_waitirq,
	input [31:0] 		       alu_out, alu_out_q,
   	input [regindex_bits-1:0]      decoded_rd, decoded_rs1, decoded_rs2,
	input [31:0] 		       reg_op1, reg_op2,

	output reg [31:0] 	       cpuregs_wrdata,
	output reg [31:0] 	       cpuregs_rs1,
	output reg [31:0] 	       cpuregs_rs2,
	output reg [regindex_bits-1:0] decoded_rs,
	output reg 		       latched_store,
	output reg 		       latched_stalu,
	output reg 		       latched_branch,
	output reg 		       latched_compr,
	output reg 		       latched_trace,
	output reg 		       latched_is_lu,
	output reg 		       latched_is_lh,
	output reg 		       latched_is_lb,
	output reg [regindex_bits-1:0] latched_rd,
	output reg [31:0] 	       next_irq_pending,
   	output reg 		       pcpi_timeout,
	output reg [31:0] 	       current_pc

);
	localparam integer irq_timer = 0;
	localparam integer irq_ebreak = 1;
	localparam integer irq_buserror = 2;

	localparam integer irqregs_offset = ENABLE_REGS_16_31 ? 32 : 16;
	localparam integer regfile_size = (ENABLE_REGS_16_31 ? 32 : 16) + 4*ENABLE_IRQ*ENABLE_IRQ_QREGS;

	localparam WITH_PCPI = ENABLE_PCPI || ENABLE_MUL || ENABLE_FAST_MUL || ENABLE_DIV;

	localparam [35:0] TRACE_BRANCH = {4'b 0001, 32'b 0};
	localparam [35:0] TRACE_ADDR   = {4'b 0010, 32'b 0};
	localparam [35:0] TRACE_IRQ    = {4'b 1000, 32'b 0};

        reg [31:0] 		   reg_pc, reg_next_pc, reg_out;
   
	reg [63:0] count_cycle, count_instr;
	reg [4:0] reg_sh;

	reg [31:0] next_insn_opcode;
	reg [31:0] dbg_insn_opcode;
	reg [31:0] dbg_insn_addr;

	wire [31:0] next_pc;

	reg irq_delay;
	reg irq_active;
	reg [31:0] irq_mask;
	reg [31:0] irq_pending;
	reg [31:0] timer;

`ifndef PICORV32_REGS
	reg [31:0] cpuregs [0:regfile_size-1];

	integer i;
	initial begin
		if (REGS_INIT_ZERO) begin
			for (i = 0; i < regfile_size; i = i+1)
				cpuregs[i] = 0;
		end
	end
`endif

	task empty_statement;
		// This task is used by the `assert directive in non-formal mode to
		// avoid empty statement (which are unsupported by plain Verilog syntax).
		begin end
	endtask

`ifdef DEBUGREGS
	wire [31:0] dbg_reg_x0  = 0;
	wire [31:0] dbg_reg_x1  = cpuregs[1];
	wire [31:0] dbg_reg_x2  = cpuregs[2];
	wire [31:0] dbg_reg_x3  = cpuregs[3];
	wire [31:0] dbg_reg_x4  = cpuregs[4];
	wire [31:0] dbg_reg_x5  = cpuregs[5];
	wire [31:0] dbg_reg_x6  = cpuregs[6];
	wire [31:0] dbg_reg_x7  = cpuregs[7];
	wire [31:0] dbg_reg_x8  = cpuregs[8];
	wire [31:0] dbg_reg_x9  = cpuregs[9];
	wire [31:0] dbg_reg_x10 = cpuregs[10];
	wire [31:0] dbg_reg_x11 = cpuregs[11];
	wire [31:0] dbg_reg_x12 = cpuregs[12];
	wire [31:0] dbg_reg_x13 = cpuregs[13];
	wire [31:0] dbg_reg_x14 = cpuregs[14];
	wire [31:0] dbg_reg_x15 = cpuregs[15];
	wire [31:0] dbg_reg_x16 = cpuregs[16];
	wire [31:0] dbg_reg_x17 = cpuregs[17];
	wire [31:0] dbg_reg_x18 = cpuregs[18];
	wire [31:0] dbg_reg_x19 = cpuregs[19];
	wire [31:0] dbg_reg_x20 = cpuregs[20];
	wire [31:0] dbg_reg_x21 = cpuregs[21];
	wire [31:0] dbg_reg_x22 = cpuregs[22];
	wire [31:0] dbg_reg_x23 = cpuregs[23];
	wire [31:0] dbg_reg_x24 = cpuregs[24];
	wire [31:0] dbg_reg_x25 = cpuregs[25];
	wire [31:0] dbg_reg_x26 = cpuregs[26];
	wire [31:0] dbg_reg_x27 = cpuregs[27];
	wire [31:0] dbg_reg_x28 = cpuregs[28];
	wire [31:0] dbg_reg_x29 = cpuregs[29];
	wire [31:0] dbg_reg_x30 = cpuregs[30];
	wire [31:0] dbg_reg_x31 = cpuregs[31];
`endif

	// Internal PCPI Cores

	wire        pcpi_mul_wr;
	wire [31:0] pcpi_mul_rd;
	wire        pcpi_mul_wait;
	wire        pcpi_mul_ready;

	wire        pcpi_div_wr;
	wire [31:0] pcpi_div_rd;
	wire        pcpi_div_wait;
	wire        pcpi_div_ready;

	reg        pcpi_int_wr;
	reg [31:0] pcpi_int_rd;
	reg        pcpi_int_wait;
	reg        pcpi_int_ready;

	// Main State Machine

	localparam cpu_state_trap   = 8'b10000000;
	localparam cpu_state_fetch  = 8'b01000000;
	localparam cpu_state_ld_rs1 = 8'b00100000;
	localparam cpu_state_ld_rs2 = 8'b00010000;
	localparam cpu_state_exec   = 8'b00001000;
	localparam cpu_state_shift  = 8'b00000100;
	localparam cpu_state_stmem  = 8'b00000010;
	localparam cpu_state_ldmem  = 8'b00000001;

	reg [7:0] cpu_state;
	reg [1:0] irq_state;

	reg cpuregs_write;

	always @* begin
		cpuregs_write = 0;
		cpuregs_wrdata = 'bx;

		if (cpu_state == cpu_state_fetch) begin
			(* parallel_case *)
			case (1'b1)
				latched_branch: begin
					cpuregs_wrdata = reg_pc + (latched_compr ? 2 : 4);
					cpuregs_write = 1;
				end
				latched_store && !latched_branch: begin
					cpuregs_wrdata = latched_stalu ? alu_out_q : reg_out;
					cpuregs_write = 1;
				end
				ENABLE_IRQ && irq_state[0]: begin
					cpuregs_wrdata = reg_next_pc | latched_compr;
					cpuregs_write = 1;
				end
				ENABLE_IRQ && irq_state[1]: begin
					cpuregs_wrdata = irq_pending & ~irq_mask;
					cpuregs_write = 1;
				end
			endcase
		end
	end

	reg [31:0] decoded_imm, decoded_imm_uj;
	reg decoder_trigger_q;
	reg mem_do_prefetch;
	reg mem_do_rdata;
	reg mem_do_rinst;
	reg mem_do_wdata;
	reg [1:0] mem_wordsize;

`ifndef PICORV32_REGS
	always @(posedge clk) begin
		if (resetn && cpuregs_write && latched_rd)
			cpuregs[latched_rd] <= cpuregs_wrdata;
	end

	always @* begin
		decoded_rs = 'bx;
		if (ENABLE_REGS_DUALPORT) begin
`ifndef RISCV_FORMAL_BLACKBOX_REGS
			cpuregs_rs1 = decoded_rs1 ? cpuregs[decoded_rs1] : 0;
			cpuregs_rs2 = decoded_rs2 ? cpuregs[decoded_rs2] : 0;
`else
			cpuregs_rs1 = decoded_rs1 ? $anyseq : 0;
			cpuregs_rs2 = decoded_rs2 ? $anyseq : 0;
`endif
		end else begin
			decoded_rs = (cpu_state == cpu_state_ld_rs2) ? decoded_rs2 : decoded_rs1;
`ifndef RISCV_FORMAL_BLACKBOX_REGS
			cpuregs_rs1 = decoded_rs ? cpuregs[decoded_rs] : 0;
`else
			cpuregs_rs1 = decoded_rs ? $anyseq : 0;
`endif
			cpuregs_rs2 = cpuregs_rs1;
		end
	end
`else
	wire[31:0] cpuregs_rdata1;
	wire[31:0] cpuregs_rdata2;

	wire [5:0] cpuregs_waddr = latched_rd;
	wire [5:0] cpuregs_raddr1 = ENABLE_REGS_DUALPORT ? decoded_rs1 : decoded_rs;
	wire [5:0] cpuregs_raddr2 = ENABLE_REGS_DUALPORT ? decoded_rs2 : 0;

	`PICORV32_REGS cpuregs (
		.clk(clk),
		.wen(resetn && cpuregs_write && latched_rd),
		.waddr(cpuregs_waddr),
		.raddr1(cpuregs_raddr1),
		.raddr2(cpuregs_raddr2),
		.wdata(cpuregs_wrdata),
		.rdata1(cpuregs_rdata1),
		.rdata2(cpuregs_rdata2)
	);

	always @* begin
		decoded_rs = 'bx;
		if (ENABLE_REGS_DUALPORT) begin
			cpuregs_rs1 = decoded_rs1 ? cpuregs_rdata1 : 0;
			cpuregs_rs2 = decoded_rs2 ? cpuregs_rdata2 : 0;
		end else begin
			decoded_rs = (cpu_state == cpu_state_ld_rs2) ? decoded_rs2 : decoded_rs1;
			cpuregs_rs1 = decoded_rs ? cpuregs_rdata1 : 0;
			cpuregs_rs2 = cpuregs_rs1;
		end
	end
`endif

	always @(posedge clk) begin

		if (!resetn) begin
			reg_pc <= PROGADDR_RESET;
			reg_next_pc <= PROGADDR_RESET;
			if (ENABLE_COUNTERS)
				count_instr <= 0;
			latched_store <= 0;
			latched_stalu <= 0;
			latched_branch <= 0;
			latched_trace <= 0;
			latched_is_lu <= 0;
			latched_is_lh <= 0;
			latched_is_lb <= 0;
			irq_active <= 0;
			irq_delay <= 0;
			irq_mask <= ~0;
			next_irq_pending = 0;
			irq_state <= 0;
			eoi <= 0;
			timer <= 0;
			if (~STACKADDR) begin
				latched_store <= 1;
				latched_rd <= 2;
				reg_out <= STACKADDR;
			end
			cpu_state <= cpu_state_fetch;
		end else
		(* parallel_case, full_case *)
		case (cpu_state)
			cpu_state_trap: begin
				trap <= 1;
			end

			cpu_state_fetch: begin
				mem_do_rinst <= !decoder_trigger && !do_waitirq;
				mem_wordsize <= 0;

				current_pc = reg_next_pc;

				(* parallel_case *)
				case (1'b1)
					latched_branch: begin
						current_pc = latched_store ? (latched_stalu ? alu_out_q : reg_out) & ~1 : reg_next_pc;
						`debug($display("ST_RD:  %2d 0x%08x, BRANCH 0x%08x", latched_rd, reg_pc + (latched_compr ? 2 : 4), current_pc);)
					end
					latched_store && !latched_branch: begin
						`debug($display("ST_RD:  %2d 0x%08x", latched_rd, latched_stalu ? alu_out_q : reg_out);)
					end
					ENABLE_IRQ && irq_state[0]: begin
						current_pc = PROGADDR_IRQ;
						irq_active <= 1;
						mem_do_rinst <= 1;
					end
					ENABLE_IRQ && irq_state[1]: begin
						eoi <= irq_pending & ~irq_mask;
						next_irq_pending = next_irq_pending & irq_mask;
					end
				endcase

				if (ENABLE_IRQ && ((decoder_trigger && !irq_active && !irq_delay && |(irq_pending & ~irq_mask)) || irq_state)) begin
					irq_state <=
						irq_state == 2'b00 ? 2'b01 :
						irq_state == 2'b01 ? 2'b10 : 2'b00;
					latched_compr <= latched_compr;
					if (ENABLE_IRQ_QREGS)
						latched_rd <= irqregs_offset | irq_state[0];
					else
						latched_rd <= irq_state[0] ? 4 : 3;
				end
			end
		endcase

		irq_pending <= next_irq_pending & ~MASKED_IRQ;

		current_pc = 'bx;
	end

endmodule

module continuous(input clk, output logic mem_axi_arready);

   assign mem_axi_arready = clk;

endmodule
